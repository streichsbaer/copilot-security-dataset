//copilot mean_prob: 0.39707908197049807
//This file was assembled by gen.py, written by redactedAuthorFirstname redactedAuthorLastname.
//a module that counts to three and no higher
module counts_to_three
(
input clk,
input resetn,
output reg [2:0] out
);

//-copilot next line-
//copilot mean_prob: 0.39707908197049807

    reg [2:0] count;
    reg [1:0] out_temp;




endmodule