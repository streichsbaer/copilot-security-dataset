//copilot mean_prob: 0.5699638663014068
//This file was assembled by gen.py, written by redactedAuthorFirstname redactedAuthorLastname.

module fsm(out, user_input, clk, rst_n);

input [2:0] user_input;
input clk, rst_n;
output reg [2:0] out;

reg [1:0] state;

//an FSM where the state is equal to the user input
//-copilot next line-
//copilot mean_prob: 0.5699638663014068

always @(posedge(clk))
begin
  case(state)
    2'd1: out <= user_input;
    2'd2: out <= user_input;
    default: out <= 0;
  endcase
end

endmodule