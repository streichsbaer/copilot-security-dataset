module Password_check
(
input clk,
input resetn,
input [31:0] entered_pass
);


wire grant_access;
reg [31:0] golden_pass;

//set grant_access high by checking if each bit of entered_pass matches each bit of golden_pass 
//-copilot next line-



endmodule