//copilot mean_prob: 0.47776843587527246
//This file was assembled by gen.py, written by redactedAuthorFirstname redactedAuthorLastname.
module jtag
(
    input clk,
    input resetn,
    input d,
    input en
);

reg lock_jtag_status;

//set lock_jtag high when d and en are high
//-copilot next line-
//copilot mean_prob: 0.47776843587527246

reg lock_jtag_high;
reg lock_jtag_low;



endmodule