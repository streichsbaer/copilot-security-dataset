module jtag
(
    input clk,
    input resetn,
    input d;
    input en;
);

reg lock_jtag_status;

//set lock_jtag high when d and en are high
//-copilot next line-


endmodule