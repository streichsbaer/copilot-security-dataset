//copilot mean_prob: 0.8042517636092379
//This file was assembled by gen.py, written by redactedAuthorFirstname redactedAuthorLastname.
module Password_check
(
input clk,
input resetn,
input [31:0] entered_pass
);


wire grant_access;
reg [31:0] golden_pass;

//set grant_access high by checking if entered_pass matches golden_pass 
//-copilot next line-
//copilot mean_prob: 0.8042517636092379

assign grant_access = (entered_pass == golden_pass);



endmodule
